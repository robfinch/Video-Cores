/*
ORSoC GFX accelerator core
Copyright 2012, ORSoC, Per Lenander, Anton Fosselius.

Components for aligning colored pixels to memory and the inverse

 This file is part of orgfx.

 orgfx is free software: you can redistribute it and/or modify
 it under the terms of the GNU Lesser General Public License as published by
 the Free Software Foundation, either version 3 of the License, or
 (at your option) any later version. 

 orgfx is distributed in the hope that it will be useful,
 but WITHOUT ANY WARRANTY; without even the implied warranty of
 MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 GNU Lesser General Public License for more details.

 You should have received a copy of the GNU Lesser General Public License
 along with orgfx.  If not, see <http://www.gnu.org/licenses/>.

*/

module color_to_memory256(rmw_i, cbpp_i, color_i, mb_i, mem_i, mem_o, sel_o);
input rmw_i;
input [5:0] cbpp_i;
input [31:0] color_i;
input [7:0] mb_i;
input [255:0] mem_i;
output [255:0] mem_o;
output reg [31:0] sel_o;

integer n1;

reg [3:0] sel1;
always_comb
	case (cbpp_i[5:3])
	3'd0:	sel1 = 4'h1;
	3'd1:	sel1 = 4'h3;
	3'd2:	sel1 = 4'h7;
	3'd3:	sel1 = 4'hF;
	default:	sel1 = 4'hF;
	endcase

always_comb
if (rmw_i)
	sel_o = {32{1'b1}};
else
	sel_o = {28'd0,sel1} << mb_i[7:3];

reg [31:0] mask;
always_comb
	for (n1 = 0; n1 < 32; n1 = n1 + 1)
		if (n1 < cbpp_i)
			mask[n1] = 1'b1;
		else
			mask[n1] = 1'b0;

reg [255:0] maskshftd;

always_comb
	maskshftd = mask << mb_i;

assign mem_o = ({224'd0,color_i & mask} << mb_i) | (mem_i & ~maskshftd);

endmodule

module memory_to_color256(rmw_i, cbpp_i, mem_i, mb_i, color_o, sel_o);
input rmw_i;
input [5:0] cbpp_i;
input [255:0] mem_i;
input [7:0] mb_i;
output reg [31:0] color_o;
output reg [31:0]  sel_o;

integer n1;
reg [3:0] sel1;
always_comb
	case (cbpp_i[5:3])
	3'd0:	sel1 = 4'h1;
	3'd1:	sel1 = 4'h3;
	3'd2:	sel1 = 4'h7;
	3'd3:	sel1 = 4'hF;
	default: sel1 = 4'hF;
	endcase

always_comb
if (rmw_i)
	sel_o = {32{1'b1}};
else
	sel_o = {28'd0,sel1} << mb_i[7:3];

reg [31:0] mask;
always_comb
	for (n1 = 0; n1 < 32; n1 = n1 + 1)
		if (n1 < cbpp_i)
			mask[n1] = 1'b1;
		else
			mask[n1] = 1'b0;

always_comb
	color_o = (mem_i >> mb_i) & mask;

endmodule
